*AM RF modulator
.AC DEC 16 1 1.0MEG
.TRAN 4U 3M
.DC VG2	LIN 1 0 10M
.PLOT V(3)
Vcc 1 0 30
VG2 2 0 DC 0 AC 1 0 SIN( 0 10M 200K 0 0 -90 )
VG1 4 0 DC 0 AC 1 0 SIN( 0 5 1K 0 0 -90 )
C3 5 0 100N
C2 6 3 470P
C1 2 7 100N
R5 0 7 15K
R4 7 1 56K
R3 0 3 1K
R2 4 5 4.7K
R1 1 6 10K
QT1 6 7 5 Q_BC548_N 
.MODEL Q_BC548_N NPN( IS=16.9F NF=1 NR=1 RE=567M RC=1
+ RB=10 VAF=56.7 VAR=28.3 ISE=154F ISC=154F 
+ NE=1.5 NC=1.5 BF=1.16K BR=5 IKF=29.5M 
+ IKR=29.5M CJC=3.35P CJE=6.85P VJC=3.57 VJE=1.09 
+ MJC=489M MJE=432M TF=796P TR=103N EG=1.11 
+ KF=0 AF=1 )
.OPTION list
.END